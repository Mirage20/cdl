

KO KOT ENF ENT ENS CN KC

ST SM

SUPF SUPC SUPT SUPCON SUPV SUPO

CLC