
Cell stock-options {
    Component stock {
        Image:Docker = "docker.io/wso2vick/sampleapp-stock"
        Ports {
             TCP 80->8080    # This is a line comment after syntax
        }
    }

    Ingress:HTTP {
        "/stock" -> stock {
            GET "/"
        }
    }
}
